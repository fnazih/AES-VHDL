    Mac OS X            	   2  �     �                                      ATTR      �     �                       com.apple.lastuseddate#PS      0   H  com.apple.macl     x  	  7com.apple.metadata:kMDLabel_y4h5lcq3l7ovlsz5rzkc6qo454     �   <  com.apple.quarantine ���]    N�     D�"�,H�>�(���                                                      ��y�ML��IHniN�L�c|Me�f�#N�
���Xjv��Ո0��/X�CE��:�C�hQ�!d4��Y�iᥟC�]�L��l������Z�"�`���U|��,�U�L�#̄�7��T����m<a��1,�-��k��/kv��L�#qϗ��#��Y�fC��A|��Ѕy���z�� V1���F��A�u�q�:�jov�*v�L
��0"ޕl��5���!���ݻa��if�	)�DvV���Y�.HdX�$>��q/0083;5dd3d301;Safari;3ABAABB0-533C-48C2-A3A8-1D2CA0985111 